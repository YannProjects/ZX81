----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09.11.2019 22:56:50
-- Design Name: 
-- Module Name: ULA - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 27-11-2021: Merge vid state machine et ULA
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use work.ZX81_Pack.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
library UNISIM;
use UNISIM.VComponents.all;
use work.ZX81_Pack.all;

entity ULA is
    Port ( CLK_3_25_M : in std_logic;
           -- Separation bus addresse CPU et RAM/ROM
           A_cpu : in std_logic_vector (15 downto 0); -- CPU address bus to ULA. Input from ULA side
           A_vid_pattern : out std_logic_vector (15 downto 0); -- Address bus to RAM/ROM memories. Output from ULA side
           -- Separation bus donnees RAM/ROM           
           D_cpu_IN : out STD_LOGIC_VECTOR (7 downto 0); -- CPU data bus IN. Output from ULA side
           D_ram_out : in STD_LOGIC_VECTOR (7 downto 0); -- RAM output data bus. Input for ULA side
           D_rom_out : in STD_LOGIC_VECTOR (7 downto 0); -- ROM ouput data bus. Input for ULA side
           -- Adresse et data vid�o pour le controlleur VGA
           vga_addr : out std_logic_vector(12 downto 0);
           vga_data : out std_logic_vector(7 downto 0);
           vga_wr_cyc : out STD_LOGIC;
           -- 
           KBDn : in STD_LOGIC_VECTOR (4 downto 0);
           TAPE_IN : in STD_LOGIC;
           USA_UK : in STD_LOGIC;
           TAPE_OUT : out STD_LOGIC;
           Iorq_Heart_Beat : out std_logic; -- Heart beat pour la sortie video
           RDn : in STD_LOGIC;
           WRn : in STD_LOGIC;
           HALTn : in STD_LOGIC;
           IORQn : in STD_LOGIC;
           NMIn : out STD_LOGIC;
           MREQn : in STD_LOGIC;
           RFRSHn : in std_logic;
           VID_PATTERN_ROM_ADDR_SELECT : out std_logic;
           M1n : in STD_LOGIC;
           WAITn : out std_logic;
           RESETn : in STD_LOGIC
         );
end ULA;

architecture Behavioral of ULA is

    type sm_video_state is (video_sm_reset, wait_for_video_exec, wait_for_m1_rfrsh, wait_for_vid_data);
    
    signal i_hsyncn : std_logic;
    signal i_vsync  : std_logic;
    signal i_nmionn : std_logic;
    signal char_line_cntr : unsigned(2 downto 0);
    signal i_vsync_pulse_duration : unsigned(11 downto 0);
    signal char_reg, vga_line_cntr, vga_line_start_offset, vga_line_start_offset_current, i_vga_data : std_logic_vector(7 downto 0);
    
    signal i_nop_detect, i_halt_detect: std_logic; 
    signal i_vga_char_offset, i_vga_addr, i_vga_rfrsh_addr : std_logic_vector(12 downto 0);
    signal i_vga_wr : std_logic;
    
    signal iorqn_0, iorqn_1, i_nmin : std_logic;
    signal i_wr_rfrsh, i_vga_rfrsh_cs : std_logic;
    
    signal state_m : sm_video_state;
    signal vid_pattern : std_logic_vector(7 downto 0);
    signal i_rom_addr_enable_for_vid_pattern, i_vsync_pulse_valid : std_logic;
    
    type sm_vga_screen_rfsh is (wait_for_screen_rfrsh_needed, rfrsh_screen_step_1, rfrsh_screen_step_2);
    signal screen_rfrsh_state_m : sm_vga_screen_rfsh;
    signal vga_line_offset_update_needed : std_logic;
    
    -- attribute mark_debug : string;
    -- attribute mark_debug of i_vsync : signal is "true";
    -- attribute mark_debug of i_vsync_pulse_valid : signal is "true";
    -- attribute mark_debug of i_hsyncn : signal is "true";
    -- attribute mark_debug of vga_addr : signal is "true";
    -- attribute mark_debug of vga_data : signal is "true";
    -- attribute mark_debug of vga_wr_cyc : signal is "true";
    -- attribute mark_debug of vga_line_start_offset : signal is "true";
   
begin

---------------------------------------------------------------------
-- Process pour la g�n�ration du HSYNC et de la gate vid�o
-- Aussi, g�n�ration du compteur de lignes par rapport au debut de la trame
---------------------------------------------------------------------
hsync_and_gate_process: process (CLK_3_25_M, RESETn)

variable hsyncn_counter: unsigned(7 downto 0);
 
begin
    if (RESETn = '0' or i_vsync = '1') then
        hsyncn_counter := X"00";
        if RESETn = '0' or i_vsync_pulse_valid = '1' then
             vga_line_cntr <= (others => '0');
        end if;
        char_line_cntr <= (others => '0');
        i_hsyncn <= '1';
    -- Sur chaque front descendant de l'horloge 6.5 MHz
    elsif rising_edge(CLK_3_25_M) then
        -- 384 cycles d'horloge � 6.5 MHz = 59 �s
        -- Duree pulse HSYNC = (414 - 384) @6.5 MHz = 4,6 �s 
        -- Generateur de HSYNC
        hsyncn_counter := hsyncn_counter + 1;
        case hsyncn_counter is
            -- HSYNCn ON 
            when FB_PORCH_OFF_DURATION =>
                i_hsyncn <= '0';
                char_line_cntr <= char_line_cntr + 1;
                vga_line_cntr <= vga_line_cntr + 1;           
            -- HSYNCn OFF
            when FB_PORCH_OFF_DURATION + HSYNC_PULSE_ON_DURATION =>
                i_hsyncn <= '1';
                hsyncn_counter := X"00";
            when others =>
                null;
        end case;
    end if;
end process;
   
-- Nouvelle version utilisant des fonctions combinatoires pour
-- le d�codage des adresses.
p_cpu_data_in : process (A_cpu, RDn, MREQn, IORQn, D_ram_out, D_rom_out, TAPE_IN, USA_UK, KBDn)
begin
    if (MREQn = '0' and RDn = '0') then
        -- Cycle de lecture RAM / ROM
        case A_cpu(15 downto 14) is
            -- Adressage de la ROM
            when "00" =>
                D_cpu_IN <= D_rom_out;
            -- Adressage de la RAM 
            when "01" =>
                D_cpu_IN <= D_ram_out;
            -- NOP execution ?
            when "11" =>
                -- NOP uniquement si le bit 6 = 0 (sinon c'est une instruction de HALT et on la laisse passer)
                if D_ram_out(6) = '0' then
                    D_cpu_IN <= X"00";
                else
                    D_cpu_IN <= D_ram_out;
                end if;
            when others =>
                D_cpu_IN <= D_rom_out;
        end case;
    elsif (IORQn = '0' and A_cpu(0) = '0' and RDn = '0') then
        -- IO inputs
        D_cpu_in <= TAPE_IN & USA_UK & '0' & KBDn(0) & KBDn(1) & KBDn(2) & KBDn(3) & KBDn(4);
    else
        D_cpu_in <= (others => 'X');
    end if;
end process;

-- Detection NOP =>  on stockera le pattern video sera lu dans la ROM dans la RAM VGA
i_nop_detect <= '1' when (M1n = '0' and MREQn = '0' and RDn = '0' and HALTn = '1' and A_cpu(15 downto 14) = "11" and D_ram_out(6) = '0') else '0';
-- Detection HALT => on stockera 0 dans la RAM VGA
i_halt_detect <= '1' when (M1n = '0' and MREQn = '0' and RDn = '0' and A_cpu(15 downto 14) = "11" and (HALTn = '0' or D_ram_out(6) = '1')) else '0';

----------------------------------------
-- Process combinatoire pour la g�n�ration ed NIMONn et VSYNC
----------------------------------------
-- Bas� sur le sch�ma http://quix.us/timex/rigter/ZX97lite.html
-- Chapitre 6) VSYNC / NMI CIRCUIT
-------------------------------------------------------
-- D'apres le schema du ZX81 clone:
-- IORQ read et A0 = 0 et NMI_ONn = 1 => VSYNC = 1
-- IORQ write => VSYNC = 0
-- IORQ write et A0 = 0 => NMI_ONn = 0 (OUT_FEn)
-- IORQ write et A1 = 0 => NMI_ONn = 1 (OUT_FDn)
-- Par rapport <E0> VSYNCn:
--          OUT_FEn => On interdit de mettre VSYNC = 1
--          OUT_FDn => On autorise de mettre VSYNC = 1
-------------------------------------------------------

-- Set/Reset pour VSYNC
p_vsync : process(RESETn, CLK_3_25_M)
begin
    if RESETn = '0' then
        i_vsync <= '0';
    -- On synchronise quand m�me avec l'horloge poursuivre les conseils de vivado 
    elsif rising_edge(CLK_3_25_M) then
        -- Enable VSYNC (IN FE)
        if IORQn = '0' and A_cpu(0) = '0' and RDn = '0' and i_nmionn = '1' then
            i_vsync <= '1';
        -- Clear VSYNC (OUT NN)
        elsif IORQn = '0' and WRn = '0' then
            i_vsync <= '0';
        end if;
    end if;    
end process;

p_vsync_pulse_duration_counter : process(RESETn, CLK_3_25_M)
begin
    if RESETn = '0' or i_vsync = '0' then
        i_vsync_pulse_duration <= X"000";
        i_vsync_pulse_valid <= '0';
    -- On compte la dur�e du pulse de VSYNC pour savoir si c'est uyne vraie synchro trame ou pas 
    elsif rising_edge(CLK_3_25_M) then
        i_vsync_pulse_duration <= i_vsync_pulse_duration + 1;
        if i_vsync_pulse_duration >= MIN_VSYNC_PULSE_DURATION then
            i_vsync_pulse_valid <= '1';
        end if;
    end if;
end process;

p_nmi : process(RESETn, CLK_3_25_M)
begin
    if RESETn = '0' then
        i_nmionn <= '1';
    -- On synchronise quand m�me avec l'horloge poursuivre les conseils de vivado        
    elsif rising_edge(CLK_3_25_M) then        
        -- Clear NMIn (OUT FD)
        if IORQn = '0' and WRn = '0' and A_cpu(1) = '0' then
            i_nmionn <= '1';
        -- Enable NMIn (OUT FE)
        elsif IORQn = '0' and WRn = '0' and A_cpu(0) = '0' then
            i_nmionn <= '0';
        end if;
    end if;
end process;

-- Process pour le comptage des caracteres par rapport au debut de la ligne 
p_vga_char_counter : process(RESETn, CLK_3_25_M, i_hsyncn)
begin
    if (RESETn = '0' or i_hsyncn = '0') then
        i_vga_char_offset <= (others => '0');
    -- Sur chaque front montant de l'horloge 3.25 MHz
    elsif rising_edge(CLK_3_25_M) then
        -- On tient compte des caracteres a afficher et aussi des instructions HALT
        -- dans ce cas, on remplira la RAM avec des 0. 
        if i_nop_detect = '1' or i_halt_detect = '1' then
            -- Incrementation de la position du caractere dans la RAM
            i_vga_char_offset <= i_vga_char_offset + 1;
        end if;
    end if;
end process;


-----------------------------------------------------
-- Process pour le heart beat IORQn (allumage LED)
-----------------------------------------------------
p_iorq_hb : process (RESETn, CLK_3_25_M, IORQn)

variable iorq_counter : unsigned(15 downto 0);
variable i_iorq_heart_beat : std_logic;

begin
    if (RESETn = '0') then
        i_iorq_heart_beat := '0';
        iorq_counter := IORQ_PERIOD;
        iorqn_1 <= '1';
    -- Sur chaque front descendant de l'horloge 6.5 MHz
    elsif rising_edge(CLK_3_25_M) then
        iorqn_0 <= IORQn;
        iorqn_1 <= iorqn_0;
        -- IORQ heart beat qui inclut le VSYNC et aussi les lectures clavier + load cassette
        -- Compteur de heart beat pour faire clignoter la LED sur le CMOD S7. 
        -- D�tection transtion 1 -> 0
        if iorqn_1 = '1' and iorqn_0 = '0' then
            iorq_counter := iorq_counter - 1;
            if  iorq_counter(15) = '1' then
                iorq_counter := IORQ_PERIOD;
                i_iorq_heart_beat := not i_iorq_heart_beat;
            end if;
        end if;
    end if;
    
    iorq_heart_beat <= i_iorq_heart_beat;
    
end process;

p_clear_screen : process  (RESETn, CLK_3_25_M, vga_line_start_offset)
begin
    if RESETn = '0' then
        screen_rfrsh_state_m <= wait_for_screen_rfrsh_needed;
        vga_line_start_offset_current <= (others => '0');
    elsif rising_edge(CLK_3_25_M) then
        case  screen_rfrsh_state_m is
            when wait_for_screen_rfrsh_needed =>
                i_vga_rfrsh_addr <= '1' & X"DFF";
                if (vga_line_start_offset /= vga_line_start_offset_current) then
                    screen_rfrsh_state_m <= rfrsh_screen_step_1;
                end if;
            when rfrsh_screen_step_1 =>
                if i_vsync_pulse_valid = '1' then
                    i_wr_rfrsh <= '1';
                    screen_rfrsh_state_m <= rfrsh_screen_step_2;
                end if;
            when rfrsh_screen_step_2 =>
                if i_vga_rfrsh_addr = X"00" then
                    vga_line_start_offset_current <= vga_line_start_offset;
                    screen_rfrsh_state_m <= wait_for_screen_rfrsh_needed;
                else
                    i_vga_rfrsh_addr <= i_vga_rfrsh_addr - 1;
                    screen_rfrsh_state_m <= rfrsh_screen_step_1;
                end if;
                i_wr_rfrsh <= '0';
            when others =>
                screen_rfrsh_state_m <= wait_for_screen_rfrsh_needed;
        end case;
    end if;
end process;
        

video_state_machine_process: process (CLK_3_25_M, RESETn)

begin
        if RESETn = '0' then
            state_m <= video_sm_reset;
        -- Sur chaque front descendant de l'horloge 6.5 MHz
        elsif rising_edge(CLK_3_25_M) then
            case state_m is
                    when video_sm_reset =>
                        i_rom_addr_enable_for_vid_pattern <= '0';
                        vga_line_start_offset <= (others => '0');
                        vga_line_offset_update_needed <= '0';
                        state_m <= wait_for_video_exec;

                     when wait_for_video_exec =>
                        i_rom_addr_enable_for_vid_pattern <= '0';
                        i_vga_wr <= '0';
                        -- Char reg contient le caract�re � afficher pr�sent dans la RAM vid�o.
                        -- Invalide en cas de HALT mais non utilis� (cas i_rom_addr_enable_for_vid_pattern = 0)
                        char_reg <= D_ram_out;
                        
                        if i_vsync = '1' and i_vsync_pulse_valid = '1' then
                             vga_line_offset_update_needed <= '1';
                        end if;

                        -- Detection front montant i_nop_detect
                        if i_nop_detect = '1' then
                            state_m <= wait_for_m1_rfrsh;
                        -- Si c'est un HALT, pas besoin de lire le pattern dans la ROM
                        elsif i_halt_detect = '1' then
                            state_m <= wait_for_vid_data;
                        end if;
                        
                     when wait_for_m1_rfrsh =>
                        if vga_line_offset_update_needed = '1' then
                            vga_line_offset_update_needed <= '0';
                            vga_line_start_offset <= vga_line_cntr;
                        end if;                  
                     
                        if RFRSHn = '0' then
                            -- Si c'est un cycle de NOP, on lit le pattern video � partir de la ROM
                            -- en construisant l'adresse � partir du caract�re � afficher et du numero
                            -- de ligne en cours.
                            A_vid_pattern <= A_cpu(15 downto 9) & char_reg(5 downto 0) & std_logic_vector(char_line_cntr(2 downto 0));
                            i_rom_addr_enable_for_vid_pattern <= '1';
                            state_m <= wait_for_vid_data;
                        end if;
                           
                     when wait_for_vid_data =>
                        if vga_line_offset_update_needed = '1' then
                            vga_line_offset_update_needed <= '0';
                            vga_line_start_offset <= vga_line_cntr;
                        end if;     
                                          
                        -- Lecture pattern vid�o
                        if i_rom_addr_enable_for_vid_pattern = '1' then
                            -- Caractere en inversion video ?
                            if (char_reg(7) = '0') then
                                vid_pattern <= D_rom_out;
                            else
                                vid_pattern <= not D_rom_out;
                            end if;
                        else
                            -- Si le CPU est en HALT, on remplit l'adresse en RAM VGA avec des 0
                            vid_pattern <= (others => '0');
                        end if;
                        
                        -- Signaux pour le controlleur VGA
                        -- Sur la totalite de la ligne, il y a 34 caract�res en tenant compte de la detection
                        -- de l'interruption de find de ligne (A_cpu(6) = 0)
                        -- Comme la RAM ne contient que 32 caract�res par ligne, on , n'ecrit pas les 2 dernier
                        -- caracteres 
                        -- if i_vga_char_offset <= 32 and vga_line_cntr > VGA_LINE_START and vga_line_cntr < VGA_LINE_STOP then
                        -- if i_vga_char_offset <= 32 and (vga_line_cntr - vga_line_start_offset >= 0)  and 
                        --     vga_line_cntr - vga_line_start_offset <= 192 then
                        if i_vga_char_offset <= 32 then
                            i_vga_wr <= '1';
                        end if;
                        state_m <= wait_for_video_exec;
                        
                     when others =>
                        state_m <= wait_for_video_exec;
            end case;
        end if;
end process;

-- Signal utilise pour postionner l'adresse du pattern video � lire en ROM
VID_PATTERN_ROM_ADDR_SELECT <= i_rom_addr_enable_for_vid_pattern;

-- Adresse de l'octet courant dans la RAM VGA. L'adresse est resette sur chaque VSYNC et incrementee quand on retourne un "NOP" ou un "HALT" au Z80
-- Adresse VGA = char_line_cntr * 32 (34 caracteres par ligne mais 32 pris en compte)  + offset caractere
i_vga_addr <= std_logic_vector(vga_line_cntr + VGA_SCREEN_OFFSET) & "00000" + i_vga_char_offset - X"1";
-- Pattern � afficher � l'ecran lu dans la ROM
i_vga_data <= vid_pattern;

vga_addr <= i_vga_rfrsh_addr when i_vga_rfrsh_cs = '1' else i_vga_addr;
vga_data <= X"00" when i_vga_rfrsh_cs = '1' else vid_pattern;
vga_wr_cyc <= i_wr_rfrsh when i_vga_rfrsh_cs = '1' else i_vga_wr;

i_vga_rfrsh_cs <= '1' when i_vsync_pulse_valid = '1' else '0';

TAPE_OUT <= not i_vsync;

-- Explications issue de la page http://www.user.dccnet.com/wrigter/index_files/ZX81WAIT.htm
-- En slow mode, le Z80 est interrompu toutes les 64 us par la NMI. La proc�dure d'interruption (en 0x0066)
-- compte le nombre de lignes restantes pour commencer l'afficahge vid�o.
-- Lorsque le nombre de ligne est atteint, le CPU ex�cute une instruction HALT et attend la prochaine NMI
-- Lorsque celle-ci arrive, le CPU continue son ex�cution � l'adresse 0x007A. Ce code, stoppe la NMI (OUT FD, A)
-- et d�mare "l'ex�cution" en RAM vid�o (JP (IX)).
-- Cependant, cette phase a besoin d'�tre synchonis�e avec la fin du pulse de NMI afin de d�marrer l'envoi
-- de la vid�o pr�ci�sement � ce moment.
-- C'est la fonction de la porte OR ci-dessous.
-- Si on sort de HALTn et que NMIn = 0 (NMI pulse en court), on ins�re des cycles de WAIT afin d'attendre la fin du pulse de NMI
-- et relacher le CPU sur le cycle T3 (apr�s les cycles de WAIT) et charger le registre � d�calage vid�o sur le cycle T4 juste apr�s...
i_nmin <= i_nmionn or i_hsyncn;
NMIn <= i_nmin;
WAITn <= not HALTn or i_nmin;

end Behavioral;
