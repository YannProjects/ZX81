----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09.11.2019 22:56:50
-- Design Name: 
-- Module Name: ULA - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 27-11-2021: Merge vid state machine et ULA
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use work.ZX81_Pack.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
library UNISIM;
use UNISIM.VComponents.all;
use work.ZX81_Pack.all;

entity ULA is
    Port ( 
           CLK_3_25_M : in std_logic;
           CLK_6_5_M : in std_logic;
           CLK_13_M : in std_logic;
           -- Separation bus addresse CPU et RAM/ROM
           A_cpu : in std_logic_vector (15 downto 0); -- CPU address bus to ULA. Input from ULA side
           A_vid_pattern : out std_logic_vector (15 downto 0); -- Address bus to RAM/ROM memories. Output from ULA side
           -- Separation bus donnees RAM/ROM           
           D_cpu_IN : out STD_LOGIC_VECTOR (7 downto 0); -- CPU data bus IN. Output from ULA side
           D_ram_out : in STD_LOGIC_VECTOR (7 downto 0); -- RAM output data bus. Input for ULA side
           D_rom_out : in STD_LOGIC_VECTOR (7 downto 0); -- ROM ouput data bus. Input for ULA side
           -- Adresse et data vid�o pour le controlleur VGA
           vga_addr : out std_logic_vector(19 downto 0);
           vga_data : out std_logic;
           vga_wr_cyc : out STD_LOGIC;
           -- 
           KBDn : in STD_LOGIC_VECTOR (4 downto 0);
           TAPE_IN : in STD_LOGIC;
           USA_UK : in STD_LOGIC;
           TAPE_OUT : out STD_LOGIC;
           vsync_heart_beat : out std_logic; -- Heart beat pour la sortie video
           RDn : in STD_LOGIC;
           WRn : in STD_LOGIC;
           HALTn : in STD_LOGIC;
           IORQn : in STD_LOGIC;
           NMIn : out STD_LOGIC;
           MREQn : in STD_LOGIC;
           RFRSHn : in std_logic;
           VID_PATTERN_ROM_ADDR_SELECT : out std_logic;
           M1n : in STD_LOGIC;
           WAITn : out std_logic;
           RESETn : in STD_LOGIC
         );
end ULA;

architecture Behavioral of ULA is

    signal i_hsyncn : std_logic;
    signal i_vsync, i_vsync_pulse_valid : std_logic;
    signal i_nmionn : std_logic;
    signal char_line_cntr : unsigned(2 downto 0);
    signal i_vsync_pulse_duration : integer;
    signal char_reg, i_d_cpu_in : std_logic_vector(7 downto 0);
    signal i_nop_detect, i_nop_detect_0: std_logic;
     
    signal i_vga_addr_frame_offset, i_vga_pixel_offset, i_vga_line_offset  : integer;
    signal i_vga_wr : std_logic;
    
    signal i_vsync_0, i_vsync_1, i_nmin : std_logic;
    
    signal i_sample_pattern_video_done : std_logic;
    
    signal i_hsyncn_cnt : integer;
    signal i_vid_shift_register : std_logic_vector(15 downto 0);
    signal i_rom_addr_enable_for_vid_pattern : std_logic;
           
    -- attribute mark_debug : string;
    -- attribute mark_debug of i_vsync : signal is "true";
    -- attribute mark_debug of i_vsync_pulse_valid : signal is "true";
    -- attribute mark_debug of i_hsyncn : signal is "true";
    -- attribute mark_debug of CLK_3_25_M : signal is "true";
    -- attribute mark_debug of CLK_6_5_M : signal is "true";
    -- attribute mark_debug of A_cpu : signal is "true";
    -- attribute mark_debug of D_cpu_IN : signal is "true";
    -- attribute mark_debug of M1n : signal is "true";
    -- attribute mark_debug of MREQn : signal is "true";
    -- attribute mark_debug of RFRSHn : signal is "true";
    -- attribute mark_debug of RDn : signal is "true";
    -- attribute mark_debug of char_line_cntr : signal is "true";
    -- attribute mark_debug of HALTn : signal is "true";
    -- attribute mark_debug of NMIn : signal is "true";
    -- attribute mark_debug of i_nmionn : signal is "true";
    -- attribute mark_debug of i_nop_detect : signal is "true";
    -- attribute mark_debug of vga_addr : signal is "true";
    -- attribute mark_debug of i_vga_addr_frame_offset : signal is "true";
    -- attribute mark_debug of i_vga_pixel_offset : signal is "true";
    -- attribute mark_debug of i_vga_line_offset : signal is "true";
    -- attribute mark_debug of vga_data : signal is "true";
    -- attribute mark_debug of vga_wr_cyc : signal is "true";

begin

p_vid_shift_register: process (CLK_13_M, RESETn)
begin
    if RESETn = '0' then
        i_vid_shift_register <= (others => '0');
        i_vga_line_offset <= 0;
    elsif rising_edge(CLK_13_M) then
        -- S�lection de la partie avec MREQn = 0 (cycle T4) durant laquelle il faut recharger le pattern video
        -- Dans le schema original du ZX81, le registre � decalage est recharge en fin de cycle T4 de l'execution en RAM video.
        -- C'est ce qui est reproduit ici en rechargeant le registre en fin de cycle T4 avec les conditions:
        -- MREQn = '0' and CLK_3_25_M = '0' and CLK_6_5_M = '0'
        -- (sur le front montant de l'horloge 13 MHz). 
        if MREQn = '0' and CLK_3_25_M = '0' and CLK_6_5_M = '0' and i_rom_addr_enable_for_vid_pattern = '1' then
            -- On resette la variable utilis�e pour adress�e une ligne ou celle du dessous avec la m�me valeur.
            i_vga_line_offset <= 0;
            -- Caractere en inversion video ?
            if (char_reg(7) = '0') then
                -- Les pixels sont doubl�s car on les �crit 2 fois:
                -- 1 fois � l'adresse A pendant le 1er cycle � 13 MHz et l'autre fois � l'adresse A + NUMBER_OF_PIXELS_PER_LINE (= nombre de pixels dans une ligne)
                -- lors du second cycle de 13 MHz. Cette solution permet de doubler les lignes verticalement.
                i_vid_shift_register <= i_d_cpu_in(7) & i_d_cpu_in(7) &
                                        i_d_cpu_in(6) & i_d_cpu_in(6) &
                                        i_d_cpu_in(5) & i_d_cpu_in(5) &
                                        i_d_cpu_in(4) & i_d_cpu_in(4) &
                                        i_d_cpu_in(3) & i_d_cpu_in(3) &
                                        i_d_cpu_in(2) & i_d_cpu_in(2) &
                                        i_d_cpu_in(1) & i_d_cpu_in(1) &
                                        i_d_cpu_in(0) & i_d_cpu_in(0) ;
            else
                i_vid_shift_register <= not (i_d_cpu_in(7) & i_d_cpu_in(7) &
                                        i_d_cpu_in(6) & i_d_cpu_in(6) &
                                        i_d_cpu_in(5) & i_d_cpu_in(5) &
                                        i_d_cpu_in(4) & i_d_cpu_in(4) &
                                        i_d_cpu_in(3) & i_d_cpu_in(3) &
                                        i_d_cpu_in(2) & i_d_cpu_in(2) &
                                        i_d_cpu_in(1) & i_d_cpu_in(1) &
                                        i_d_cpu_in(0) & i_d_cpu_in(0)) ;
            end if;
        else
            if i_vga_line_offset = 0 then
                -- Ligne du dessous (1 cycle de 13 MHz sur 2)
                i_vga_line_offset <= NUMBER_OF_PIXELS_PER_LINE;
            else
                -- Ligne courante (1 cycle de 13 MHz sur 2)
                i_vga_line_offset <= 0;
            end if;
            i_vid_shift_register <= i_vid_shift_register(14 downto 0) & '0';
        end if;
    end if;
end process;

p_vga_addr_counter: process (CLK_6_5_M, i_vsync, RESETn)
begin
    if RESETn = '0' or i_hsyncn = '0' or i_vsync = '1' then
        -- On resette le nombre de pixel depuis le d�but de la ligne en cas de HSYNCn ou VSYNC
        i_vga_pixel_offset <= 0;
    elsif rising_edge(CLK_6_5_M) then
        -- On d�bute le comptage des pixels  de ligne a partir du moment ou on a atteind
        -- la fin du pulse de VSYNC
        if i_hsyncn_cnt < FB_PORCH_OFF_DURATION then
            -- On incremente de 2 pixels pour doubler le nombre de pixels de ligne
            i_vga_pixel_offset <= i_vga_pixel_offset + 2;
        end if;
    end if;
end process;

-- i_vga_addr_frame_offset: Adresse du d�but de la la ligne courante dans la trame
-- i_vga_pixel_offset: Offset du pixel dans la ligne
-- i_vga_line_offset: Variable utilis�e pour adress�e un ligne sur 2 (contient 0 ou NUMBER_OF_PIXELS_PER_LINE)
-- LINE_OFFSET_FROM_FRAME_START: Offset pour d�caler l'image de 45 lignes vers le haut et mieux la centrer par rapport � l'affichage VGA
-- PIXEL_LINE_START: Offset dans la ligne du premier pixel � �crire
-- PIXEL_LINE_STOP: Offset dans la ligne du dernier pixel � �crire
-- Une ligne d'affichage du ZX81 contient 192 cycles d'horloge � 3,5 MHz donc 384 cycles � 6,5 MHz, soit un maximum de 384 pixels par lignes.
-- Si on double l'affichage pour utiliser la totalit� de la ligne de 640x480, on arrive � 384 * 2 > 640 pixels, 
-- le mieux est d'�liminer les premiers et dernier pixels pour n'avoir que 640 pixels par ligne:
-- 2*384 - 640 = 128. J'ai donc mis 64 PIXEL_LINE_START ce qui correspond � 64 pixels de ligne VGA sur la partie gauche qui sont elimines de la ligne.

vga_addr <= std_logic_vector(to_unsigned(i_vga_addr_frame_offset + i_vga_pixel_offset + i_vga_line_offset - FRAME_LINE_START - PIXEL_LINE_START, vga_addr'length));
vga_data <= i_vid_shift_register(15);
vga_wr_cyc <= i_hsyncn and not i_vsync when i_vga_addr_frame_offset >= FRAME_LINE_START and 
                                            i_vga_pixel_offset >= PIXEL_LINE_START and
                                            i_vga_pixel_offset < PIXEL_LINE_STOP 
                                       else '0';

---------------------------------------------------------------------
-- Process pour la g�n�ration du HSYNC et de la gate vid�o
-- Aussi, g�n�ration du compteur de lignes par rapport au debut de la trame
---------------------------------------------------------------------
hsync_and_gate_process: process (CLK_3_25_M, RESETn)

variable hsyncn_counter: integer;
 
begin
    if (RESETn = '0' or i_vsync = '1') then
        hsyncn_counter := 0;
        char_line_cntr <= (others => '0');
        if (RESETn = '0' or i_vsync_pulse_valid = '1') then
            i_vga_addr_frame_offset <= 0;
        end if;
        i_hsyncn <= '1';
    -- Sur chaque front descendant de l'horloge 3,25 MHz
    elsif rising_edge(CLK_3_25_M) then
        -- 192 cycles d'horloge � 3,25 MHz
        -- Duree pulse HSYNC = (207 - 192) @3,25 MHz = 4,6 �s 
        hsyncn_counter := hsyncn_counter + 1;
        if hsyncn_counter >= FB_PORCH_OFF_DURATION and hsyncn_counter < FB_PORCH_OFF_DURATION + HSYNC_PULSE_ON_DURATION then  
            i_hsyncn <= '0';
        elsif hsyncn_counter = FB_PORCH_OFF_DURATION + HSYNC_PULSE_ON_DURATION then
            i_hsyncn <= '1';
            char_line_cntr <= char_line_cntr + 1;
            i_vga_addr_frame_offset <= i_vga_addr_frame_offset + 2*NUMBER_OF_PIXELS_PER_LINE;
            hsyncn_counter := 0;
        end if;
    end if;
    
    i_hsyncn_cnt <= hsyncn_counter;
    
end process;

-- Nouvelle version utilisant des fonctions combinatoires pour
-- le d�codage des adresses.
p_cpu_data_in : process (A_cpu, RDn, MREQn, IORQn, RFRSHn, D_ram_out, D_rom_out, TAPE_IN, USA_UK, KBDn)
begin
    -- MREQn = '0' and RFRSHn = '0' pour tenir compte du mode HiRers o� l'on doit pouvoir lire des patterns
    -- video � partir de la RAM et pas seulement de la ROM.
    if (MREQn = '0' and RDn = '0') or (MREQn = '0' and RFRSHn = '0') then
        -- Cycle de lecture RAM / ROM
        case A_cpu(15 downto 14) is
            -- Adressage de la ROM
            when "00" =>
                i_d_cpu_in <= D_rom_out;
            -- Adressage de la RAM 
            when "01" =>
                i_d_cpu_in <= D_ram_out;
            -- NOP execution ?
            when "11" =>
                -- NOP uniquement si le bit 6 = 0 (sinon c'est une instruction de HALT et on la laisse passer)
                if D_ram_out(6) = '0' then
                    i_d_cpu_in <= X"00";
                else
                    i_d_cpu_in <= D_ram_out;
                end if;
            when others =>
                i_d_cpu_in <= D_rom_out;
        end case;
    elsif (IORQn = '0' and A_cpu(0) = '0' and RDn = '0') then
        -- IO inputs
        i_d_cpu_in <= TAPE_IN & USA_UK & '0' & KBDn(0) & KBDn(1) & KBDn(2) & KBDn(3) & KBDn(4);
    else
        i_d_cpu_in <= (others => 'X');
    end if;
end process;

D_cpu_in <= i_d_cpu_in;

-- Detection NOP =>  on stockera le pattern video sera lu dans la ROM dans la RAM VGA
i_nop_detect <= '1' when (M1n = '0' and MREQn = '0' and RDn = '0' and HALTn = '1' and A_cpu(15 downto 14) = "11" and D_ram_out(6) = '0') else '0';

----------------------------------------
-- Process combinatoire pour la g�n�ration ed NIMONn et VSYNC
----------------------------------------
-- Bas� sur le sch�ma http://quix.us/timex/rigter/ZX97lite.html
-- Chapitre 6) VSYNC / NMI CIRCUIT
-------------------------------------------------------
-- D'apres le schema du ZX81 clone:
-- IORQ read et A0 = 0 et NMI_ONn = 1 => VSYNC = 1
-- IORQ write => VSYNC = 0
-- IORQ write et A0 = 0 => NMI_ONn = 0 (OUT_FEn)
-- IORQ write et A1 = 0 => NMI_ONn = 1 (OUT_FDn)
-- Par rapport <E0> VSYNCn:
--          OUT_FEn => On interdit de mettre VSYNC = 1
--          OUT_FDn => On autorise de mettre VSYNC = 1
-------------------------------------------------------

-- Set/Reset pour VSYNC
p_vsync : process(RESETn, CLK_3_25_M)
begin
    if RESETn = '0' then
        i_vsync <= '0';
    -- On synchronise quand m�me avec l'horloge poursuivre les conseils de vivado 
    elsif rising_edge(CLK_3_25_M) then
        -- Enable VSYNC (IN FE)
        if IORQn = '0' and A_cpu(0) = '0' and RDn = '0' and i_nmionn = '1' then
            i_vsync <= '1';
        -- Clear VSYNC (OUT NN)
        elsif IORQn = '0' and WRn = '0' then
            i_vsync <= '0';
        end if;
    end if;    
end process;

p_vsync_pulse_duration_counter : process(RESETn, CLK_3_25_M)
begin
    if RESETn = '0' or i_vsync = '0' then
        i_vsync_pulse_duration <= 0;
        i_vsync_pulse_valid <= '0';
    -- On compte la dur�e du pulse de VSYNC pour savoir si c'est uyne vraie synchro trame ou pas
    -- (cas du ZX81 en mode pseudo-hires avec invaders ou pacman)
    elsif rising_edge(CLK_3_25_M) then
        i_vsync_pulse_duration <= i_vsync_pulse_duration + 1;
        if i_vsync_pulse_duration >= MIN_VSYNC_PULSE_DURATION then
            i_vsync_pulse_valid <= '1';
        end if;
    end if;
end process;

p_nmi : process(RESETn, CLK_3_25_M)
begin
    if RESETn = '0' then
        i_nmionn <= '1';
    -- On synchronise quand m�me avec l'horloge poursuivre les conseils de vivado        
    elsif rising_edge(CLK_3_25_M) then        
        -- Clear NMIn (OUT FD)
        if IORQn = '0' and WRn = '0' and A_cpu(1) = '0' then
            i_nmionn <= '1';
        -- Enable NMIn (OUT FE)
        elsif IORQn = '0' and WRn = '0' and A_cpu(0) = '0' then
            i_nmionn <= '0';
        end if;
    end if;
end process;

-----------------------------------------------------
-- Process pour le heart beat (allumage LED)
-----------------------------------------------------
p_vsync_hb : process (RESETn, CLK_3_25_M, IORQn)

variable i_vsync_counter : integer;
variable i_heart_beat : std_logic;

begin
    if (RESETn = '0') then
        i_heart_beat := '0';
        i_vsync_counter := VSYNC_COUNTER_PERIOD;
    -- Sur chaque front descendant de l'horloge 6.5 MHz
    elsif rising_edge(CLK_3_25_M) then
        i_vsync_0 <= i_vsync_pulse_valid;
        i_vsync_1 <= i_vsync_0;
        -- Compteur de heart beat pour faire clignoter la LED sur le CMOD S7. 
        -- D�tection transtion 1 -> 0
        if i_vsync_1 = '1' and i_vsync_0 = '0' then
            i_vsync_counter := i_vsync_counter - 1;
            if  i_vsync_counter = 0 then
                i_vsync_counter := VSYNC_COUNTER_PERIOD;
                i_heart_beat := not i_heart_beat;
            end if;
        end if;
    end if;
    
    vsync_heart_beat <= i_heart_beat;
    
end process;
        
nop_detect_process: process (CLK_3_25_M)
begin
    if rising_edge(CLK_3_25_M) then
        -- Le signalde NOP est d�cal� de 2 p�riodes de 3,25 MHz
        -- pour se caler sur les cycles CPU T3 et T4
        i_nop_detect_0 <= i_nop_detect;
        -- Le signal est align� sur les cycle T3 et T4 de l'execution en RAM pour l'affichage video
        i_rom_addr_enable_for_vid_pattern <= i_nop_detect_0;
        -- Si NOP detect, on lit le caract�re dans la RAM
        if i_nop_detect = '1' then
            char_reg <= D_ram_out;
        end if;
    end if;
end process;

A_vid_pattern <= A_cpu(15 downto 9) & char_reg(5 downto 0) & std_logic_vector(char_line_cntr);
-- Signal utilise pour positionner l'adresse du pattern video � lire en ROM
VID_PATTERN_ROM_ADDR_SELECT <= i_rom_addr_enable_for_vid_pattern;

TAPE_OUT <= not i_vsync;

-- Explications issue de la page https://quix.us/timex/rigter/ZX97lite.html
-- En slow mode, le Z80 est interrompu toutes les 64 us par la NMI. La proc�dure d'interruption (en 0x0066)
-- compte le nombre de lignes restantes pour commencer l'affichage vid�o.
-- Lorsque le nombre de ligne est atteint, le CPU ex�cute une instruction HALT et attend la prochaine NMI
-- Lorsque celle-ci arrive, le CPU continue son ex�cution � l'adresse 0x007A. Ce code, stoppe la NMI (OUT FD, A)
-- et d�mare "l'ex�cution" en RAM vid�o (JP (IX)).
-- Cependant, cette phase a besoin d'�tre synchonis�e avec la fin du pulse de NMI afin de d�marrer l'envoi
-- de la vid�o pr�ci�sement � ce moment.
-- C'est la fonction de la porte OR ci-dessous.
-- Si on sort de HALTn et que NMIn = 0 (NMI pulse en court), on ins�re des cycles de WAIT afin d'attendre la fin du pulse de NMI
-- et relacher le CPU sur le cycle T3 (apr�s les cycles de WAIT) et charger le registre � d�calage vid�o sur le cycle T4 juste apr�s...
i_nmin <= i_nmionn or i_hsyncn;
NMIn <= i_nmin;
WAITn <= not HALTn or i_nmin;

end Behavioral;
