----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09.11.2019 22:56:50
-- Design Name: 
-- Module Name: ULA - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 27-11-2021: Merge vid state machine et ULA
-- 02-04-2023: Redesign the ULA to be closer to ZX97 (https://quix.us/timex/rigter/ZX97lite.html)
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use work.ZX81_Pack.all;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
library UNISIM;
use UNISIM.VComponents.all;
use work.ZX81_Pack.all;

entity ULA is
    Port ( 
           i_resetn : in std_logic;
           
           -- System clocks
           i_clk_3_25_m : in std_logic;
           i_clk_6_5_m : in std_logic;
           
           i_A : in std_logic_vector(15 downto 0);
           
           -- A'[8..0] addresses generated by ULA
           o_Ap : out std_logic_vector(8 downto 0);
           
           -- Character index inside ZX81 RAM or pattern data inside ZX81 ROM
           i_video_pattern : in std_logic_vector(7 downto 0);
           
           -- ULA data (NOP or I/O: KBD, Tape in,...)
           o_ula_data : out std_logic_vector(7 downto 0);
           
           -- Keyboard raws
           i_kbdn : in std_logic_vector (4 downto 0);
           
           -- Load/Save
           i_tape_in : in std_logic;
           i_usa_uk : in std_logic;
           o_tape_out : out std_logic;

           o_ram_csn : out std_logic;
           o_rom_csn : out std_logic;
           -- Put ULA data to Z80
           o_ulan : out std_logic;
           
           -- Z80 control signals
           i_rdn : in std_logic;
           i_wrn : in std_logic;
           i_haltn : in std_logic;
           i_iorqn : in std_logic;
           i_mreqn : in std_logic;
           i_m1n : in std_logic;
           i_rfshn : in std_logic;
           o_waitn : out std_logic;
           o_nmin : out std_logic;
                      
           -- Video
           o_vsync : out std_logic;
           o_hsync : out std_logic;
           o_video_data : out std_logic
           
         );
end ULA;

architecture Behavioral of ULA is

    signal hsync, hsync0, hsync1 : std_logic;
    signal vsync : std_logic;
    signal nmionn, kbd_n : std_logic;
    signal char_line_cntr : unsigned(2 downto 0);
    signal char_reg : std_logic_vector(7 downto 0);
    signal nop_detect, nmin : std_logic;
    signal reload_vid_pattern : std_logic;
     
    signal vid_shift_register : std_logic_vector(7 downto 0);
    
    signal hsyncn_counter : unsigned(7 downto 0);
    signal nop_delay : std_logic_vector(2 downto 0);
    
begin

-- U14, U13.A, U13.B, U23.C
p_memory_decoder: process (i_rdn, i_rfshn, i_mreqn, i_A, i_m1n)
begin
    if (i_rfshn and i_mreqn) = '0' then
        case i_A(15 downto 14) is
            -- 0x0000 -> 0x1FFF (8K)
            when "00" =>
                o_ram_csn <= '1';
                o_rom_csn <= '0';
            -- 0x4000 -> 0x6FFF (16K)
            -- 0xC000 -> 0xFFFF (Video memory)
            when "01"|"10" =>
                o_ram_csn <= '0';
                o_rom_csn <= '1';
            when "11" =>
                o_ram_csn <= i_m1n;
                o_rom_csn <= not i_m1n;                                 
            when others =>
                o_ram_csn <= '1';
                o_rom_csn <= '1';
        end case;
    else
        o_ram_csn <= '1';
        o_rom_csn <= '1';
    end if;
end process;

-- CHR$ decoder
-- U11
p_chr_decoder: process (i_clk_3_25_m, i_resetn, vsync)
begin
    if i_resetn = '0' or vsync = '1' then
        char_line_cntr <= (others => '0');
    elsif rising_edge(i_clk_3_25_m) then
        hsync1 <= hsync;
        hsync0 <= hsync1;
        -- HSYNC falling edge 
        if hsync0 = '1' and hsync1 = '0' then
            char_line_cntr <= char_line_cntr + 1;
        end if;
    end if;
end process;

-- U12
o_Ap <= char_reg(5 downto 0) & std_logic_vector(char_line_cntr) when i_rdn = '0';

-- Timing generator
p_hsync_gen: process (i_clk_3_25_m, i_resetn, vsync)
begin
    -- 192 cycles d'horloge � 3,25 MHz
    if i_resetn = '0' or vsync = '1' or hsyncn_counter = FB_PORCH_OFF_DURATION + HSYNC_PULSE_ON_DURATION then
        hsyncn_counter <= X"00";
    elsif rising_edge(i_clk_3_25_m) then
        hsyncn_counter <= hsyncn_counter + 1;
    end if;
end process;

-- Duree pulse HSYNC = (207 - 192) @3,25 MHz = 4,6 �s 
hsync <= '1' when hsyncn_counter >= FB_PORCH_OFF_DURATION else '0';

----------------------------------------
-- Process combinatoire pour la g�n�ration ed NIMONn et VSYNC
----------------------------------------
-- Bas� sur le sch�ma http://quix.us/timex/rigter/ZX97lite.html
-- Chapitre 6) VSYNC / NMI CIRCUIT
-------------------------------------------------------
-- D'apres le schema du ZX97:
-- IORQ read et A0 = 0 et NMI_ONn = 1 => VSYNC = 1
-- IORQ write => VSYNC = 0
-- IORQ write et A0 = 0 => NMI_ONn = 0 (OUT_FEn)
-- IORQ write et A1 = 0 => NMI_ONn = 1 (OUT_FDn)
-- Par rapport <E0> VSYNCn:
--          OUT_FEn => On interdit de mettre VSYNC = 1
--          OUT_FDn => On autorise de mettre VSYNC = 1
-------------------------------------------------------

-- VSYNC NMI KBD (U8, U15, U17)
p_vsync : process(i_iorqn, i_A, i_rdn, i_wrn)
begin
    -- Clear VSYNC (OUT NN)
    if (i_iorqn = '0' and i_wrn = '0') or i_resetn = '0' then
        vsync <= '0';
    -- Enable VSYNC (IN FE)
    elsif i_iorqn = '0' and i_A(0) = '0' and i_rdn = '0' then
        vsync <= '1';
    end if;
end process;

p_nmi : process(i_iorqn, i_A, i_rdn, i_wrn)
begin
    -- Clear NMIn (OUT FD)
    if (i_iorqn = '0' and i_wrn = '0' and i_A(1) = '0') or i_resetn = '0' then
        nmionn <= '1';
    -- Enable NMIn (OUT FE)
    elsif i_iorqn = '0' and i_wrn = '0' and i_A(0) = '0' then
        nmionn <= '0';
    end if;
end process;

-- Explications issue de la page https://quix.us/timex/rigter/ZX97lite.html
-- En slow mode, le Z80 est interrompu toutes les 64 us par la NMI. La proc�dure d'interruption (en 0x0066)
-- compte le nombre de lignes restantes pour commencer l'affichage vid�o.
-- Lorsque le nombre de ligne est atteint, le CPU ex�cute une instruction HALT et attend la prochaine NMI
-- Lorsque celle-ci arrive, le CPU continue son ex�cution � l'adresse 0x007A. Ce code, stoppe la NMI (OUT FD, A)
-- et d�mare "l'ex�cution" en RAM vid�o (JP (IX)).
-- Cependant, cette phase a besoin d'�tre synchonis�e avec la fin du pulse de NMI afin de d�marrer l'envoi
-- de la vid�o pr�cis�ement � ce moment.
-- C'est la fonction de la porte OR ci-dessous.
-- Si on sort de HALTn et que NMIn = 0 (NMI pulse en court), on ins�re des cycles de WAIT afin d'attendre la fin du pulse de NMI
-- et relacher le CPU sur le cycle T3 (apr�s les cycles de WAIT) et charger le registre � d�calage vid�o sur le cycle T4 juste apr�s...
nmin <= nmionn or not hsync;
o_waitn <= not i_haltn or nmin;
o_nmin <= nmin;

-- Lecture entr�e clavier (U8)
kbd_n <= (i_A(0) or i_rdn) or i_iorqn;
o_ulan <= not(not kbd_n or nop_detect);
o_ula_data <= i_TAPE_IN & i_USA_UK & '0' & i_kbdn(0) & i_kbdn(1) & i_kbdn(2) & i_kbdn(3) & i_kbdn(4) when kbd_n = '0' else (others => '0');
o_tape_out <= not vsync;

-- NOP detection (U19, U13)
nop_detect <= '1' when (i_m1n = '0' and i_mreqn = '0' and i_rdn = '0' and i_haltn = '1' and i_A(15 downto 14) = "11" and i_video_pattern(6) = '0') else '0';
char_reg <= i_video_pattern when nop_detect = '1';

-- Retarde le NOP de 2 cycles de 6,5 MHz pour �tre synchonis� avec l'instant de rechargement du 
-- pattern video
p_process_nop_delay: process(i_clk_6_5_m)
begin
    if rising_edge(i_clk_6_5_m) then
        nop_delay <= nop_delay(1 downto 0) & nop_detect;
    end if;
end process;

reload_vid_pattern <= '1' when nop_delay="100" else '0';

-- Registre � d�calage (U22)
p_vid_shift_register: process (i_clk_6_5_m, reload_vid_pattern)
begin
    if rising_edge(i_clk_6_5_m) then
        if reload_vid_pattern = '1' then
            -- Caractere en inversion video ?
            if (char_reg(7) = '0') then
                vid_shift_register <= i_video_pattern;
            else
                vid_shift_register <= not i_video_pattern;
            end if;
        else
            vid_shift_register <= vid_shift_register(6 downto 0) & '0';
        end if;
    end if;
end process;

o_video_data <= vid_shift_register(7);
o_hsync <= hsync;
o_vsync <= vsync;

end Behavioral;
